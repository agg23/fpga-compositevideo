`define PLL_DYN
`define PLL_DEVICE "GW1NR-9C"
`define PLL_FCLKIN "27"
